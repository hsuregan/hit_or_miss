/*
this module is in between frequency and randomizer,
everytime frequency sends a pulse to this module,
a random number comes up
*/

